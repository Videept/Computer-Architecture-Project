module displayA
(
    input[5:0] x,
    output[5:0] y
);
//This module is to set ouptut as first 8 bit number    
assign y=x;
endmodule
